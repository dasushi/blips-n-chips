module mips(input clk, reset,
					input logic [31:0] instr_addr, instr_in, data_out,
					output logic [31:0] data_addr, data_in,
					output logic data_rd_wr); //1=read
	parameter [31:0] pc_init = 32'h80020000;
    parameter [31:0] sp_init = 32'h80120000; //= 32'h80020000 + 2**20
	parameter [31:0] ra_init = 32'h00000000;
    
	logic [4:0] instr_counter; //Rolling bit counter to detect which stage the instruction is in
	logic [31:0] mem_index; // Offset address for next block of bytes in multi word reads
	logic [31:0] pc; // corrected address removes the 8002xxxx from MIPS compiled hexadecimal
	logic [31:0] instr_reg;
	logic [31:0] mem_reg;
	
	regfile #() regs(.wr_num(), .wr_data(), wr_en(),
		.rd0_num(), .rd0_data(),
		.rd1_num(), .rd1_data(),
		.clk(clk));
	//instructions we will need: 	
	//addiu addu jr li lw move nop sw
	//pages refer to pdf page # in MIPS ISA
	
	//ADDI rt, rs, immediate
	//add immediate unsigned (pg 47)
	
	//ADDU rd, rs, rt
	//add unsigned word (pg 48)
	
	//JR rs
	//jump register, set PC to rs (pg 155)
	
	//LI rt, immediate
	//load immediate to reg (not in ISA - is this upper or lower? or full 32 bit?)
	
	//LW rt, offset(base)
	//load word to memory (pg 171)
	
	//MOVE rd, rs
	//move register to register
	
	//NOP
	//not an op, actually SLL r0, r0, 0 (pg 226)
	
	//SW, rt, offset(base)
	//store word from rt to memory[base+offset] (pg 280)
	
	initial begin
		//initialize
	end
	
	always @ ( access_size, addr, rd_wr) begin
		if(enable && rd_wr) begin
			byte_offset = addr[1:0];
			set_mem_index(addr); 
			word_counter = 4'h0;
			read_data(mem_index, byte_offset, 4'd0);
		end else begin
			if(~rd_wr) begin
				data_out = 32'bx;
			end
		end
	end
	
	//main task
	always @ (posedge clk)
	begin : STAGES
		// Determine which stage
		case(instr_counter)
			5'b00001 : begin //IF
				instr_addr <= pc;
				mem_reg <= instr_in;
				instr_reg <= mem_reg;
				pc <= pc + 32h'00000004;
			end
			5'b00010 : begin //ID
				//decode current_instr to instruction (+ immediate)
			end
			5'b00100 : begin //EX
				//execute arithmetic, eg. address = base + offset
			end
			5'b01000 : begin //ME
				//read from calculated address
			end
			5'b10000 : begin //WB
				//write back to memory if required
			end
			endcase
		end
		instr_counter <= instr_counter << 1;
	end // clock
	
	//may still be useful
	task set_mem_index(input [31:0] address);
	begin
		mem_index = addr ^ 32'h80020000; // Clear the base address generated by MIPS compiler
		mem_index = mem_index - byte_offset;
		mem_index = mem_index >> 2; // Takes the Floor (integer division) 
	end
	endtask

endmodule