module mips(input clk, reset,
					input logic [31:0] instr_addr, instr_in, data_out,
					output logic [31:0] data_addr, data_in,
					output logic data_rd_wr); //1=read
	parameter [31:0] pc_init = 32'h80020000;
    parameter [31:0] sp_init = 32'h80120000; //= 32'h80020000 + 2**20
	parameter [31:0] ra_init = 32'h00000000;
    
	logic reg_wr_en, alu_en, wb_en, mem_en;
	logic [4:0] instr_counter,	//Rolling bit counter to detect which stage the instruction is in
				wr_sel, rt_sel, rs_sel;
	logic [31:0] pc; 			// program counter
	logic [31:0] instr_reg, 	// current instruction register
				 em_reg, 		// memory data register (mdr/mbr)
				 rt, 			// register output 1
				 rs, 			// register output 2
				 rd, 			// destination register
				 alu_1, 		// alu input 1
				 alu_2, 		// alu input 2
				 alu_out,		// alu output reg
	regfile #() regs(.wr_num(wr_sel), .wr_data(rd), wr_en(reg_wr_en),
		.rd0_num(rt_sel), .rd0_data(rt),
		.rd1_num(rs_sel), .rd1_data(rs),
		.clk(clk));
	
	initial begin
		//initialize
	end
	
	//main task
	always @ (posedge clk)
	begin : STAGES
		// Determine which stage
		case(instr_counter)
			5'b00001 : begin //IF
				instr_addr <= pc;
				mem_reg <= instr_in;
				instr_reg <= mem_reg;
				pc <= pc + 32h'00000004;
			end
			5'b00010 : begin //ID
				//decode current_instr to instruction (+ immediate)
				//instructions we will need: 	
				//addiu addu jr li lw move nop sw
				//pages refer to pdf page # in MIPS ISA
				case(instr_reg[31:26])
					6b'001001 : begin //ADDIU
					//ADDIU rt, rs, immediate
					//add immediate unsigned (pg 47)
					//[31:26]: 001001
					wr_sel <= instr_reg[20:16]; //store result here (rt)
					rs_sel <= instr_reg[25:21]; //operand 1, rs 
					alu_1 <= rs;
					sign_extend(instr_reg[15:0]); //operand 2, immediate, sets alu_2
					alu_en <= 1'b1;
					wb_en <= 1'b1;
					end
					
					6b'100011 : begin //LW
					//LW rt, offset(base)
					//load word to memory (pg 171) 
					//[31:26]: 100011
					wr_sel <= instr_reg[20:16]; // store from mem to this reg (rt)
					rd_sel <= instr_reg[25:21]; // base addr
					alu_1 <= rd;
					sign_extend(instr_reg[15:0]); //sets alu_2 with offset
					alu_en <= 1'b1;
					end
					
					//NOTE: LW and SW seem similar so far - change to common stage? only diff is 10(0/1)011
					6b'101011 : begin //SW
					//SW, rt, offset(base)
					//store word from rt to memory[base+offset] (pg 280)
					//address error exception if last two bits != 00
					//[31:26]: 101011
					rt_sel <= instr_reg[20:16]; //source word
					rd_sel <= instr_reg[25:21]; //base address
					alu_1 <= rd;
					sign_extend(instr_reg[15:0]); //sets alu_2 with immediate
					alu_en <= 1'b1;
					end
					
					6b'000000 : begin //SPECIAL
					case(instr_reg[5:0]) 
						6'b100001 : begin //ADDU
						//ADDU rd, rs, rt
						//add unsigned word (pg 48)
						//[31:26]: 000000 & [5:0]: 100001
						rs_sel <= instr_reg[25:21];
						rt_sel <= instr_reg[20:16];
						rd_sel <= instr_reg[15:11];
						end
						6'b001000 : begin
						//JR rs
						//jump register, set PC to rs (pg 155) 
						//[31:26]: 000000 & [5:0]: 0010000
						end
						6'b001000 : begin
						//LI rt, immediate
						//load immediate to reg (not in ISA - is this upper or lower? or full 32 bit?)
						end
						6'b001000 : begin
						//MOVE rd, rs
						//move register to register
						end
						6'b000000 : begin
						//NOP
						//not an op, actually SLL r0, r0, 0 (pg 226) do we need to actually implement this way?
						//[31:26]: 000000 & SLL [5:0]=000000
						end
					end
				end
			end
			5'b00100 : begin //EX
				//execute arithmetic and instruction, eg. address = base + offset
				//run if alu_en is set
				//adds alu_1 and alu_2
				//output to alu_out
				if(alu_en == 1'b1) begin
					alu_out <= alu_1 + alu_2;
				end
			end
			5'b01000 : begin //ME
				//read from calculated address
			end
			5'b10000 : begin //WB
				//write back to memory if required
			end
			endcase
		end
		instr_counter <= instr_counter << 1;
	end // clock
	
	//may still be useful
	task set_mem_index(input [31:0] address);
	begin
		mem_index = addr ^ 32'h80020000; // Clear the base address generated by MIPS compiler
		mem_index = mem_index - byte_offset;
		mem_index = mem_index >> 2; // Takes the Floor (integer division) 
	end
	endtask
	
	task sign_extend(input [15:0] val);
	begin
		//TODO: determine what reg to write to (ALU input 2)
		alu_2[31:16] <= (val[15]===1'b1) ? 16h'ffff : 16h'0000; //sign extend with 1 if neg, 0 if pos
		alu_2[15:0] <= val;
	end
	endtask

endmodule