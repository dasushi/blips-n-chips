module memory(input clk,
					input logic [31:0] addr, data_in,
					output logic [31:0] data_out,
					input logic [1:0] access_size,
					input logic rd_wr,
					output logic busy,
					input logic enable);
	parameter benchmark = "whatever.x";
    parameter depth = 2**20; // =1 MB
    
	reg[0:31] mem [depth-1: 0];
	logic [4:0] word_counter; //Rolling bit counter to detect offest/ which word is next to be read for multi word reads
	logic [1:0] byte_offset;
	logic [31:0] mem_index; // Offset address for next block of bytes in multi word reads
	logic [31:0] base_address; // corrected address removes the 8002xxxx from MIPS compiled hexadecimal
	
	initial begin
		$readmemh(benchmark, mem);
		busy = 0;
		byte_offset = 0;
		word_counter = 5'd0;
		byte_offset = addr[1:0];
		set_mem_index(addr);
		base_address = 32'b0;
	end

	always @ (addr) begin
		byte_offset = addr[1:0];
		set_mem_index(addr); 
	end

	task set_mem_index(input [31:0] address);
	begin
		mem_index = addr ^ 32'h80020000; // Clear the base address generated by MIPS compiler
		mem_index = mem_index - byte_offset;
		mem_index = mem_index >> 2; // Takes the Floor (integer division) 
	end
	endtask
	
	always @ (posedge clk)
	begin : READ
		if(enable && rd_wr) begin
				// Read operations
				case(access_size)
					2'b00 : begin	// 4 Byte Read (Word)
						read_data(byte_offset);
					end
					2'b01 : begin	// 16 bytes (4 Words) 
						busy = 1;

						read_data(byte_offset);
						mem_index = mem_index + 1;
						word_counter = word_counter + 5'd1;
						// reset word counter if completed read
						if(word_counter == 5'd4) begin
							word_counter = 5'b0;
							busy = 0;
							set_mem_index(addr);
						end
					end
					2'b10: begin	// 32 Bytes (8 Words)
						busy = 1;

						read_data(byte_offset);

						mem_index = mem_index + 1;

						word_counter = word_counter + 5'd1;
						// reset word counter if completed read
						if(word_counter == 5'd8) begin
							word_counter = 5'b0;
							busy = 0;
							set_mem_index(addr);
						end
					end
					2'b11: begin
						// 64 Bytes (16 Words)
						busy = 1;

						read_data(byte_offset);

						mem_index = mem_index + 1;
						word_counter = word_counter + 5'd1;
						// reset word counter if completed read
						if(word_counter == 5'd16) begin
							word_counter = 5'b0;
							busy = 0;
							set_mem_index(addr);
						end
					end
					endcase
		end
	end // clock
	
	always @ (posedge clk) 
	begin : WRITE
		if(enable && ~rd_wr) begin	
			write_data(byte_offset);
		end
	end
	

	task read_data(input logic[1:0] byte_offset);
	begin
		case(byte_offset)
			2'h0: begin
				data_out = mem[mem_index];
			end
			2'h1: begin
				data_out = {mem[mem_index][8:31],  mem[mem_index + 1][0:7]};
			end
			2'h2: begin
				data_out = {mem[mem_index][16:31],  mem[mem_index+1][0:15]};
			end
			2'h3: begin
				data_out = {mem[mem_index][24:31],  mem[mem_index+1][0:23]};
			end
		endcase
	end
	endtask

	task write_data(input logic[1:0] byte_offset);
	begin
		case(byte_offset)
		2'h0: begin
			//Default Word write
			mem[mem_index] = data_in;
		end
		2'h1: begin
			mem[mem_index] = {mem[mem_index][24:31], data_in[31:8]};
			mem[mem_index + 1][24:31] = data_in[7:0];
		end
		2'h2: begin
			mem[mem_index] = {mem[mem_index][15:31], data_in[31:16]};
			mem[mem_index + 1][16:31] = data_in[15:0];
		end
		2'h3: begin
			mem[mem_index] = {mem[mem_index][0:7],data_in[31:24]};
			mem[mem_index + 1] = {mem[mem_index][8:31], data_in[23:0]};
		end
		endcase
	end
	endtask

endmodule