module memory(input clk,
					input logic [31:0] addr, data_in,
					output logic [31:0] data_out,
					input logic [1:0] access_size,
					input logic rd_wr,
					output logic busy,
					input logic enable);
	parameter benchmark = "whatever.x";
    parameter depth = 2**20; // =1 MB
    
	reg[0:31] mem [depth-1: 0];
	logic [3:0] word_counter; //Rolling bit counter to detect offest/ which word is next to be read for multi word reads
	logic [4:0] next_word_counter;
	logic [1:0] byte_offset;
	logic [31:0] mem_index; // Offset address for next block of bytes in multi word reads
	logic [31:0] base_address; // corrected address removes the 8002xxxx from MIPS compiled hexadecimal
	
	initial begin
		$readmemh(benchmark, mem);
		busy = 0;
		byte_offset = 0;
		word_counter = 5'd0;
		byte_offset = addr[1:0];
		set_mem_index(addr);
		base_address = 32'b0;
	end
	
	always @ (enable, access_size, addr, rd_wr) begin
		if(enable && rd_wr) begin
			byte_offset = addr[1:0];
			set_mem_index(addr); 
			word_counter = 4'h0;
			read_data(mem_index, byte_offset, 4'd0);
		end
	end

	task set_mem_index(input [31:0] address);
	begin
		mem_index = addr ^ 32'h80020000; // Clear the base address generated by MIPS compiler
		mem_index = mem_index - byte_offset;
		mem_index = mem_index >> 2; // Takes the Floor (integer division) 
	end
	endtask
	
	always @ (posedge clk)
	begin : READ

		if(enable && rd_wr) begin
				// Read operations
				case(access_size)
					2'b00 : begin	// 4 Byte Read (Word)
						read_data(mem_index, byte_offset, 4'h0);
						word_counter = 4'h0;
					end
					2'b01 : begin	// 16 bytes (4 Words) 
						busy = 1;
						
						read_data(mem_index, byte_offset, word_counter + 5'd1);
						word_counter = word_counter + 5'd1;

						// reset word counter if completed read
						if(word_counter == 4'h3) begin
							word_counter = 4'h0;
							busy = 0;
							set_mem_index(addr);
						end
					end
					2'b10: begin	// 32 Bytes (8 Words)
						busy = 1;

						read_data(mem_index, byte_offset, word_counter + 5'd1);
						word_counter = word_counter + 5'd1;

						// reset word counter if completed read
						if(word_counter == 4'h7) begin
							word_counter = 4'h0;
							busy = 0;
							set_mem_index(addr);
						end
					end
					2'b11: begin
						// 64 Bytes (16 Words)
						busy = 1;
					    read_data(mem_index, byte_offset, word_counter + 5'd1);
						word_counter = word_counter + 5'd1;

						// reset word counter if completed read
						if(word_counter == 4'hf) begin
							word_counter = 4'h0;
							busy = 0;
							set_mem_index(addr);
						end
					end
					endcase
		end
	end // clock
	
	always @ (posedge clk) 
	begin : WRITE
		if(enable && ~rd_wr) begin	
			write_data(byte_offset);
		end
	end
	

	task read_data(input logic [31:0] address , input logic[1:0] byte_offset, logic[3:0] word_counter);
	begin
		case(byte_offset)
			2'h0: begin
				data_out = mem[address + word_counter];
			end
			2'h1: begin
				data_out = {mem[address + word_counter][8:31],  mem[address + word_counter + 1][0:7]};
			end
			2'h2: begin
				data_out = {mem[address + word_counter][16:31],  mem[address + word_counter + 1][0:15]};
			end
			2'h3: begin
				data_out = {mem[address + word_counter][24:31],  mem[address + word_counter + 1][0:23]};
			end
		endcase
	end
	endtask

	task write_data(input logic[1:0] byte_offset);
	begin
		case(byte_offset)
		2'h0: begin
			//Default Word write
			mem[mem_index] = data_in;
		end
		2'h1: begin // Fills 1,2,3 + 4
			mem[mem_index] = {mem[mem_index][0:7],data_in[31:8]};
			mem[mem_index + 1] = {data_in[7:0], mem[mem_index][8:31]};
		end
		2'h2: begin	// Fills 2,3, + 4,5
			mem[mem_index] = {mem[mem_index][0:15],data_in[31:16]};
			mem[mem_index + 1] = {data_in[15:0], mem[mem_index][16:31]};
		end
		2'h3: begin // Fills 3 + 4,5,6
			mem[mem_index] = {mem[mem_index][0:23],data_in[31:24]};
			mem[mem_index + 1] = {data_in[23:0], mem[mem_index][24:31]};
		end
		endcase
	end
	endtask

endmodule