module mips(input clk, reset,
					input logic [31:0] instr_addr, instr_in, data_addr, data_in, 
					output logic [31:0] data_out,
					input logic data_rd_wr);
	parameter [31:0] pc_init = 32'h80020000;
    parameter [31:0] sp_init = 32'h80120000; //= 32'h80020000 + 2**20
	parameter [31:0] ra_init = 32'h00000000;
    
	logic [4:0] instr_counter; //Rolling bit counter to detect which stage the instruction is in
	logic [31:0] mem_index; // Offset address for next block of bytes in multi word reads
	logic [31:0] base_address; // corrected address removes the 8002xxxx from MIPS compiled hexadecimal
	regfile #() regs(.wr_num(), .wr_data(), wr_en(),
		.rd0_num(), .rd0_data(),
		.rd1_num(), .rd1_data(),
		.clk(clk));
		
	//addiu addu jr li lw move nop sw
	//ADDI rt, rs, immediate
	//add immediate unsigned (pg 47)
	//ADDU rd, rs, rt
	//add unsigned word (pg 48)
	//JR rs
	//jump register, set PC to rs (pg 155)
	//LI rt, immediate
	//load immediate to reg (not in ISA - is this upper or lower? or full 32 bit?)
	//LW rt, offset(base)
	//load word to memory (pg 171)
	//MOVE rd, rs
	//move register to register
	//NOP
	//not an op, actually SLL r0, r0, 0 (pg 226)
	//SW, rt, offset(base)
	//store word from rt to memory[base+offset] (pg 280)
	
	initial begin
		//initialize
	end
	
	always @ ( access_size, addr, rd_wr) begin
		if(enable && rd_wr) begin
			byte_offset = addr[1:0];
			set_mem_index(addr); 
			word_counter = 4'h0;
			read_data(mem_index, byte_offset, 4'd0);
		end else begin
			if(~rd_wr) begin
				data_out = 32'bx;
			end
		end
	end
	
	//main task
	always @ (posedge clk)
	begin : STAGES
		// Determine which stage
		case(instr_counter)
			5'b00000 : begin
			end
			5'b00001 : begin
			end
			5'b00010 : begin	
			end
			5'b00100 : begin
			end
			5'b01000 : begin
			end
			5'b10000 : begin
			end
			endcase
		end
	end // clock
	
	//may still be useful
	task set_mem_index(input [31:0] address);
	begin
		mem_index = addr ^ 32'h80020000; // Clear the base address generated by MIPS compiler
		mem_index = mem_index - byte_offset;
		mem_index = mem_index >> 2; // Takes the Floor (integer division) 
	end
	endtask

	task read_data(input logic [31:0] address , input logic[1:0] byte_offset, logic[3:0] word_counter);
	begin
		case(byte_offset)
			2'h0: begin
				data_out = mem[address + word_counter];
			end
			2'h1: begin
				data_out = {mem[address + word_counter][8:31],  mem[address + word_counter + 1][0:7]};
			end
			2'h2: begin
				data_out = {mem[address + word_counter][16:31],  mem[address + word_counter + 1][0:15]};
			end
			2'h3: begin
				data_out = {mem[address + word_counter][24:31],  mem[address + word_counter + 1][0:23]};
			end
		endcase
	end
	endtask

	task write_data(input logic[1:0] byte_offset);
	begin
		case(byte_offset)
		2'h0: begin
			//Default Word write
			mem[mem_index] = data_in;
		end
		2'h1: begin // Fills 1,2,3 + 4
			mem[mem_index] = {mem[mem_index][0:7],data_in[31:8]};
			mem[mem_index + 1] = {data_in[7:0], mem[mem_index][8:31]};
		end
		2'h2: begin	// Fills 2,3, + 4,5
			mem[mem_index] = {mem[mem_index][0:15],data_in[31:16]};
			mem[mem_index + 1] = {data_in[15:0], mem[mem_index][16:31]};
		end
		2'h3: begin // Fills 3 + 4,5,6
			mem[mem_index] = {mem[mem_index][0:23],data_in[31:24]};
			mem[mem_index + 1] = {data_in[23:0], mem[mem_index][24:31]};
		end
		endcase
	end
	endtask

endmodule